library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity DF_5to32_Decoder is
    Port ( D_IN : in STD_LOGIC_VECTOR(4 downto 0);
           F_OUT : out STD_LOGIC_VECTOR(31 downto 0);
           enable : in std_logic);
end DF_5to32_Decoder;

architecture Dataflow of DF_5to32_Decoder is

begin

    -- Dataflow modeling with 'with ... select'
    F_OUT <= "00000000000000000000000000000000" when enable = '0' else  --If enable is 0, F_OUT is set to all zeroes
             "00000000000000000000000000000001" when D_IN = "00000" else
             "00000000000000000000000000000010" when D_IN = "00001" else
             "00000000000000000000000000000100" when D_IN = "00010" else
             "00000000000000000000000000001000" when D_IN = "00011" else
             "00000000000000000000000000010000" when D_IN = "00100" else
             "00000000000000000000000000100000" when D_IN = "00101" else
             "00000000000000000000000001000000" when D_IN = "00110" else
             "00000000000000000000000010000000" when D_IN = "00111" else
             "00000000000000000000000100000000" when D_IN = "01000" else
             "00000000000000000000001000000000" when D_IN = "01001" else
             "00000000000000000000010000000000" when D_IN = "01010" else
             "00000000000000000000100000000000" when D_IN = "01011" else
             "00000000000000000001000000000000" when D_IN = "01100" else
             "00000000000000000010000000000000" when D_IN = "01101" else
             "00000000000000000100000000000000" when D_IN = "01110" else
             "00000000000000001000000000000000" when D_IN = "01111" else
             "00000000000000010000000000000000" when D_IN = "10000" else
             "00000000000000100000000000000000" when D_IN = "10001" else
             "00000000000001000000000000000000" when D_IN = "10010" else
             "00000000000010000000000000000000" when D_IN = "10011" else
             "00000000000100000000000000000000" when D_IN = "10100" else
             "00000000001000000000000000000000" when D_IN = "10101" else
             "00000000010000000000000000000000" when D_IN = "10110" else
             "00000000100000000000000000000000" when D_IN = "10111" else
             "00000001000000000000000000000000" when D_IN = "11000" else
             "00000010000000000000000000000000" when D_IN = "11001" else
             "00000100000000000000000000000000" when D_IN = "11010" else
             "00001000000000000000000000000000" when D_IN = "11011" else
             "00010000000000000000000000000000" when D_IN = "11100" else
             "00100000000000000000000000000000" when D_IN = "11101" else
             "01000000000000000000000000000000" when D_IN = "11110" else
             "10000000000000000000000000000000" when D_IN = "11111";

end Dataflow;

